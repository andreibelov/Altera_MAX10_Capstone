-- Entity
entity C4M1P1 is port (
  i_clk             : in  std_logic;
  i_data            : in  std_logic_vector(7 downto 0);
  o_parity          : out std_logic);
end entity C4M1P1;

-- Architecture
architecture rtl of C4M1P1 is begin
end architecture rtl;
